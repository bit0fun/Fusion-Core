module add(reg_a, reg_b, sum, flg_carry, flg_zero, carryin);

	parameter NBIT = 32;

	input[(NBIT-1):0] reg_a, reg_b;
	input carryin;
	output[(NBIT-1):0] sum;

	output flg_carry, flg_zero;

	wire[(NBIT-1):0] bit_sum; 	//only 1 bit, make
	wire[(NBIT-1):0] p;	    	//values for fast carry
	wire[(NBIT-1):0] g;
	wire[(NBIT):0] carry;	//intermediary carry bits
	
	/*Carry generator intermediary step*/
	wire[(NBIT):1] carry_p; 	//p[n] & p[n-1] & ... & carryin
	wire[(NBIT):1] carry_g;	//(g[0] & p[n] & p[n-1]...)


	genvar i; //for counter

	begin
	for(i = 0; i <= NBIT; i = i+1)
		assign g[i] = reg_a[i] & reg_b[i];
	end

	begin
	for(i = 0; i <= NBIT; i = i+1)
		assign p[i] = reg_a[i] | reg_b[i];
	end


	/*Intermediary Carry Assignments*/
	begin
		assign carry_p[1]  = p[0] & carryin;
		assign carry_p[2]  = p[0] & p[1] & carryin;
		assign carry_p[3]  = p[0] & p[1] & p[2] & carryin;
		assign carry_p[4]  = p[0] & p[1] & p[2] & p[3] & carryin;
		assign carry_p[5]  = p[0] & p[1] & p[2] & p[3] & p[4] & carryin;
		assign carry_p[6]  = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & carryin;
		assign carry_p[7]  = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & carryin;
		assign carry_p[8]  = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & carryin;
		assign carry_p[9]  = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & carryin;
		assign carry_p[10] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & carryin;
		assign carry_p[11] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & carryin;
		assign carry_p[12] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & carryin;
		assign carry_p[13] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & carryin;
		assign carry_p[14] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] carryin;
		assign carry_p[15] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & carryin;
		assign carry_p[16] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & carryin;
		assign carry_p[17] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & carryin;
		assign carry_p[18] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & carryin;
		assign carry_p[19] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & carryin;
		assign carry_p[20] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & carryin;
		assign carry_p[21] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12]
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & carryin;
		assign carry_p[22] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & carryin;
		assign carry_p[23] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & carryin;
		assign carry_p[24] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & carryin;
		assign carry_p[25] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] 
				 & carryin;
		assign carry_p[26] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] 
				 & p[25] & carryin;
		assign carry_p[27] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] 
				 & p[25] & p[26] & carryin;
		assign carry_p[28] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] 
				 & p[25] & p[26] & p[27] & carryin;
		assign carry_p[29] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] 
				 & p[25] & p[26] & p[27] & p[28] & carryin;
		assign carry_p[30] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] 
				 & p[25] & p[26] & p[27] & p[28] & p[29] & carryin;
		assign carry_p[31] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] 
				 & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & carryin;
		assign carry_p[32] = p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] 
				 & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] 
				 & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31] & carryin;
	end

	begin
		assign carry_g[1] = g[0];
		assign carry_g[2] = (g[0] & p[1]) + g[1];
		assign carry_g[3] = (g[0] & p[1] & p[2]) + (g[1] & p[2]) + g[2];
		assign carry_g[4] = (g[0] & p[1] & p[2] & p[3]) + (g[1] & p[2] & p[3]) + (g[2] & p[3]) + g[3];
		assign carry_g[5] = (g[0] & p[1] & p[2] & p[3] & p[4]) + (g[1] & p[2] & p[3] & p[4]) + (g[2] & p[3] & p[4]) + (g[3] & p[4]) + g[4];
		assign carry_g[6] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5]) + (g[1] & p[2] & p[3] & p[4] & p[5]) + (g[2] & p[3] & p[4] & p[5]) 
			+ (g[3] & p[4] & p[5]) + (g[4] & p[5]) + g[5];
		assign carry_g[7] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6]) + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]) + (g[2] & p[3] & p[4] & p[5] & p[6]) 
			+ (g[3] & p[4] & p[5] & p[6]) + (g[4] & p[5] & p[6]) + (g[5] & p[6]) + g[6];
		assign carry_g[8] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7]) + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7]) + (g[3] & p[4] & p[5] & p[6] & p[7]) + (g[4] & p[5] & p[6] & p[7]) 
			+ (g[5] & p[6] & p[7]) + (g[6] & p[7]) + g[7];
		assign carry_g[9] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8]) + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8]) + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8]) + (g[4] & p[5] & p[6] & p[7] & p[8]) 
			+ (g[5] & p[6] & p[7] & p[8]) + (g[6] & p[7] & p[8]) + (g[7] & p[8]) + g[8];
		assign carry_g[10] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9]) + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9]) + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9]) + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9]) + (g[6] & p[7] & p[8] & p[9]) + (g[7] & p[8] & p[9]) + (g[8] & p[9]) + g[9];
		assign carry_g[11] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10]) + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10]) + (g[6] & p[7] & p[8] & p[9] & p[10]) + (g[7] & p[8] & p[9] & p[10])
		        + (g[8] & p[9] & p[10]) + (g[9] & p[10]) + g[10];
		assign carry_g[12] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11]) + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11]) + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11])
		        + (g[7] & p[8] & p[9] & p[10]& p[11])
		        + (g[8] & p[9] & p[10] & p[11]) + (g[9] & p[10] & p[11]) + (g[10] & p[11]) + g[11];
		assign carry_g[13] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12])
		        + (g[8] & p[9] & p[10] & p[11] & p[12])
		        + (g[9] & p[10] & p[11] & p[12]) + (g[10] & p[11] & p[12]) + (g[11] & p[12]) + g[12];
		assign carry_g[14] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13])
		        + (g[9] & p[10] & p[11] & p[12] & p[13])
			+ (g[10] & p[11] & p[12] & p[13]) + (g[11] & p[12] & p[13]) + (g[12] & p[13]) + g[13];
		assign carry_g[15] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14])
			+ (g[10] & p[11] & p[12] & p[13] & p[14])
			+ (g[11] & p[12] & p[13] & p[14]) + (g[12] & p[13] & p[14]) + (g[13] & p[14]) + g[14];

		/*16 BITS FINISHED*/

		assign carry_g[16] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15])
			+ (g[11] & p[12] & p[13] & p[14] & p[15])
			+ (g[12] & p[13] & p[14] & p[15]) + (g[13] & p[14] & p[15]) + (g[14] & p[15]) + g[15];
		assign carry_g[17] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16])
			+ (g[12] & p[13] & p[14] & p[15] & p[16])
			+ (g[13] & p[14] & p[15] & p[16]) + (g[14] & p[15] & p[16]) + (g[15] & p[16]) + g[16];
		assign carry_g[18] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17])
			+ (g[13] & p[14] & p[15] & p[16] & p[17])
			+ (g[14] & p[15] & p[16] & p[17]) + (g[15] & p[16] & p[17]) + (g[16] & p[17]) + g[17];
		assign carry_g[19] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18])
			+ (g[14] & p[15] & p[16] & p[17] & p[18])
			+ (g[15] & p[16] & p[17] & p[18]) + (g[16] & p[17] & p[18]) + (g[17]  & p[18]) + g[18];
		assign carry_g[20] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19])
			+ (g[14] & p[15] & p[16] & p[17] & p[18] & p[19])
			+ (g[15] & p[16] & p[17] & p[18] & p[19])
			+ (g[16] & p[17] & p[18] & p[19]) + (g[17]  & p[18] & p[19]) + (g[18] & p[19]) + g[19];
		assign carry_g[21] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20])
			+ (g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20])
			+ (g[16] & p[17] & p[18] & p[19] & p[20])
			+ (g[17]  & p[18] & p[19] & p[20]) + (g[18] & p[19] & p[20]) + (g[19] & p[20]) + g[20];
		assign carry_g[22] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20] & p[21])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
			+ (g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21])
			+ (g[16] & p[17] & p[18] & p[19] & p[20] & p[21])
			+ (g[17]  & p[18] & p[19] & p[20] & p[21])
			+ (g[18] & p[19] & p[20] & p[21]) + (g[19] & p[20] & p[21]) + (g[20] & p[21]) + g[21];
		assign carry_g[23] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
			+ (g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
			+ (g[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22])
			+ (g[17]  & p[18] & p[19] & p[20] & p[21] & p[22])
			+ (g[18] & p[19] & p[20] & p[21] & p[22])
			+ (g[19] & p[20] & p[21] & p[22]) + (g[20] & p[21] & p[22]) + (g[21] & p[22]) + g[22];

		assign carry_g[24] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
			+ (g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
			+ (g[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
			+ (g[17]  & p[18] & p[19] & p[20] & p[21] & p[22] & p[23])
			+ (g[18] & p[19] & p[20] & p[21] & p[22] & p[23])
			+ (g[19] & p[20] & p[21] & p[22] & p[23])
			+ (g[20] & p[21] & p[22] & p[23]) + (g[21] & p[22] & p[23]) + (g[22] & p[23]) + g[23];
		assign carry_g[25] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
			+ g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
			+ (g[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
			+ (g[17]  & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
			+ (g[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24])
			+ (g[19] & p[20] & p[21] & p[22] & p[23] & p[24])
			+ (g[20] & p[21] & p[22] & p[23] & p[24])
			+ (g[21] & p[22] & p[23] & p[24]) + (g[22] & p[23] & p[24]) + (g[23] & p[24]) + g[24];

		assign carry_g[26] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[17]  & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[20] & p[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[21] & p[22] & p[23] & p[24] & p[25])
			+ (g[22] & p[23] & p[24] & p[25]) + (g[23] & p[24] & p[25]) + (g[24] & p[25]) + g[25];

		assign carry_g[27] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[17]  & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[21] & p[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[22] & p[23] & p[24] & p[25] & p[26])
			+ (g[23] & p[24] & p[25] & p[26]) + (g[24] & p[25] & p[26]) + (g[25] & p[26]) + g[26];

		assign carry_g[28] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[17]  & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[22] & p[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[23] & p[24] & p[25] & p[26] & p[27])
			+ (g[24] & p[25] & p[26] & p[27]) + (g[25] & p[26] & p[27]) + (g[26] & p[27]) + g[27];

		assign carry_g[29] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[17]  & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[23] & p[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[24] & p[25] & p[26] & p[27] & p[28])
			+ (g[25] & p[26] & p[27] & p[28]) + (g[26] & p[27] & p[28]) + (g[27] & p[28]) + g[28];

		assign carry_g[30] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[17]  & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[24] & p[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[25] & p[26] & p[27] & p[28] & p[29])
			+ (g[26] & p[27] & p[28] & p[29]) + (g[27] & p[28] & p[29]) + (g[28] & p[29]) + g[29];
		assign carry_g[31] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[17]  & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[25] & p[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[26] & p[27] & p[28] & p[29] & p[30])
			+ (g[27] & p[28] & p[29] & p[30]) + (g[28] & p[29] & p[30]) + (g[29] & p[30]) + g[30];
		assign carry_g[32] = (g[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
		        + (g[1] & p[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31]) 
			+ (g[2] & p[3] & p[4] & p[5] & p[6]& p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31]) 
		        + (g[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
		        + (g[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31]) 
			+ (g[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
		        + (g[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
		        + (g[7] & p[8] & p[9] & p[10]& p[11] & p[12] & p[13] & p[14] & p[15 & p[16]] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
		        + (g[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
		        + (g[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ g[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[17]  & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[26] & p[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[27] & p[28] & p[29] & p[30] & p[31])
			+ (g[28] & p[29] & p[30] & p[31]) + (g[29] & p[30] & p[31]) + (g[30] & p[31]) + g[31];

	end

	/*Carry assignments*/
	begin
		assign carry[0]  = carryin;
		assign carry[1]  = carry_p[1] + carry_g[1];
		assign carry[2]  = carry_p[2] + carry_g[2];
		assign carry[3]  = carry_p[3] + carry_g[3];
		assign carry[4]  = carry_p[4] + carry_g[4];
		assign carry[5]  = carry_p[5] + carry_g[5];
		assign carry[6]  = carry_p[6] + carry_g[6];
		assign carry[7]  = carry_p[7] + carry_g[7];
		assign carry[8]  = carry_p[8] + carry_g[8];
		assign carry[9]  = carry_p[9] + carry_g[9];
		assign carry[10]  = carry_p[10] + carry_g[10];
		assign carry[11]  = carry_p[11] + carry_g[11];
		assign carry[12]  = carry_p[12] + carry_g[12];
		assign carry[13]  = carry_p[13] + carry_g[13];
		assign carry[14]  = carry_p[14] + carry_g[14];
		assign carry[15]  = carry_p[15] + carry_g[15];
		assign carry[16]  = carry_p[16] + carry_g[16];
		assign carry[17]  = carry_p[17] + carry_g[17];
		assign carry[18]  = carry_p[18] + carry_g[18];
		assign carry[19]  = carry_p[19] + carry_g[19];
		assign carry[20]  = carry_p[20] + carry_g[20];
		assign carry[21]  = carry_p[21] + carry_g[21];
		assign carry[22]  = carry_p[22] + carry_g[22];
		assign carry[23]  = carry_p[23] + carry_g[23];
		assign carry[24]  = carry_p[24] + carry_g[24];
		assign carry[25]  = carry_p[25] + carry_g[25];
		assign carry[26]  = carry_p[26] + carry_g[26];
		assign carry[27]  = carry_p[27] + carry_g[27];
		assign carry[28]  = carry_p[28] + carry_g[28];
		assign carry[29]  = carry_p[29] + carry_g[29];
		assign carry[30]  = carry_p[30] + carry_g[30];
		assign carry[31]  = carry_p[31] + carry_g[31];
		assign carry[32]  = carry_p[32] + carry_g[32];
	end



always@*
	begin
	
	end



endmodule
